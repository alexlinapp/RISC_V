module aludec
    (
        input logic         opb5,
        input logic [2:0]   funct3,
        input logic         funct7b5,
        input logic [1:0]   ALUOp,
        output logic [2:0]  ALUControl
    );
    logic RTypeSub;
   
endmodule
