`include "uvm_macros.svh"
package scoreboard_pkg
    
endpackage