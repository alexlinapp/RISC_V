package global_defs_pkg;
    parameter int XLEN = 32;
    parameter int DMEM_SIZE = 64; //  max number of words memory can hold
    parameter int IMEM_SIZE = 64;
endpackage