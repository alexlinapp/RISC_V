module hazardunit
    (
        
        
        output  logic                   StallF, StallD,
        output  logic                   FlushE,
        output  logic [1:0]             ForwardAE, ForwardBE
    );
endmodule
