package callback_pkg;


    class className extends superClass;
        function new();
            
        endfunction //new()
    endclass //className extends superClass
endpackage